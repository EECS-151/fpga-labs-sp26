module one_bit_comparator_always (
    input logic a,
    input logic b,
    output logic greater,
    output logic less,
    output logic equal
);
    always_comb begin
        if (____) begin // TODO
            // TODO
        end else if (____) begin // TODO
            // TODO
        end else begin
            // TODO
        end
    end
endmodule