module one_bit_comparator_structural (
    input  logic a,
    input  logic b,
    output logic greater,
    output logic less,
    output logic equal
);
    logic a_not, b_not;

    not(____); // TODO
    not(____); // TODO

    and(________); // TODO
    and(________); // TODO
    xnor(________); // TODO
endmodule