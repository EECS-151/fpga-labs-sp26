module four_bit_comparator_always (
    input ____ a, // TODO
    input ____ b, // TODO
    output logic greater,
    output logic less,
    output logic equal
);
    always_comb begin
        if (____) begin // TODO
            // TODO
        end else if (____) begin // TODO
            // TODO
        end else begin
            // TODO
        end
    end
endmodule