module one_bit_comparator_behavioral (
    input  logic a,
    input  logic b,
    output logic greater,
    output logic less,
    output logic equal
);
    ____ greater = ________; // TODO
    ____ less    = ________; // TODO
    ____ equal   = ________; // TODO
endmodule