module edge_detector #(
    parameter WIDTH = 1
)(
    input logic clk,
    input logic [WIDTH-1:0] signal_in,
    output logic [WIDTH-1:0] edge_detect_pulse
);
    // TODO: Implement a multi-bit edge detector that detects a rising edge of 'signal_in[x]'
    // and outputs a one-cycle pulse 'edge_detect_pulse[x]' at the next clock edge
    // Feel free to use as many number of registers you like

    // Remove this line once you create your edge detector
    assign edge_detect_pulse = 0;
endmodule
