module synchronizer #(parameter int WIDTH = 1) (
    input wire [WIDTH-1:0] async_signal,
    input wire clk,
    output logic [WIDTH-1:0] sync_signal
);
    // TODO: Create your 2 flip-flop synchronizer here
    // This module takes in a vector of WIDTH-bit asynchronous
    // (from different clock domain or not clocked, such as button press) signals
    // and should output a vector of WIDTH-bit synchronous signals
    // that are synchronized to the input clk

    // Remove this line once you create your synchronizer
    assign sync_signal = 0;
endmodule
