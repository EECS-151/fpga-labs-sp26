module line_decoder (
    input  logic [3:0] select,
    input  logic [3:0] addr,
    output logic       single_wire
);
    assign single_wire = ________; // TODO
endmodule